// module mcu_fpga_bus (
    
// );
    
// endmodule